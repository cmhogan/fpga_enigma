// Copyright (c) 2026, Chad Hogan
// All rights reserved.
// Use of this source code is governed by a BSD-style
// license that can be found in the LICENSE file.

// plugboard_tb.v
// — Self-checking testbench for FPGA Enigma I plugboard commands
// Tests :S-- (plugboard clear) and re-wiring after clear
// Architecture: A continuous background UART receiver deposits bytes into
// a FIFO. The main test sequence pulls bytes via get_byte. This avoids
// send/receive timing overlap issues.

`timescale 1ns / 1ps

module plugboard_tb;

    // =========================================================================
    // Clock and DUT
    // =========================================================================
    reg clk = 1'b0;
    always #41.667 clk = ~clk;  // ~12 MHz (83.333 ns period)

    reg  uart_rx_pin = 1'b1;    // idle HIGH
    wire uart_tx_pin;
    wire led_d1, led_d2, led_d3, led_d4, led_d5;

    enigma_top dut (
        .clk       (clk),
        .ext_rst_n (1'b1),
        .uart_rx   (uart_rx_pin),
        .uart_tx   (uart_tx_pin),
        .led_d1    (led_d1),
        .led_d2    (led_d2),
        .led_d3    (led_d3),
        .led_d4    (led_d4),
        .led_d5    (led_d5)
    );

    // =========================================================================
    // VCD dump for coverage
    // =========================================================================
    `ifdef VCD_DUMP
    initial begin
        $dumpfile("build/plugboard_tb.vcd");
        $dumpvars(0, plugboard_tb);
    end
    `endif

    // =========================================================================
    // Baud rate constants
    // =========================================================================
    localparam BAUD_CLKS = 104;  // 12MHz / 115200 ≈ 104

    // =========================================================================
    // Background UART receiver → byte FIFO
    // =========================================================================
    reg [7:0] rx_fifo [0:255];
    integer   rx_wr_ptr = 0;
    integer   rx_rd_ptr = 0;

    // Continuous receiver: runs forever, depositing bytes into rx_fifo
    initial begin : bg_receiver
        reg [7:0] shift;
        integer bi;
        forever begin
            @(negedge uart_tx_pin);   // wait for start bit
            repeat(BAUD_CLKS / 2) @(posedge clk);  // midpoint of start bit
            shift = 8'd0;
            for (bi = 0; bi < 8; bi = bi + 1) begin
                repeat(BAUD_CLKS) @(posedge clk);
                shift = {uart_tx_pin, shift[7:1]};
            end
            repeat(BAUD_CLKS) @(posedge clk);  // stop bit
            rx_fifo[rx_wr_ptr[7:0]] = shift;
            rx_wr_ptr = rx_wr_ptr + 1;
        end
    end

    // get_byte: blocks until a byte is available, then returns it
    task get_byte;
        output [7:0] data;
        begin
            wait(rx_rd_ptr < rx_wr_ptr);
            data = rx_fifo[rx_rd_ptr[7:0]];
            rx_rd_ptr = rx_rd_ptr + 1;
        end
    endtask

    // =========================================================================
    // Test counters
    // =========================================================================
    integer pass_count = 0;
    integer fail_count = 0;
    integer test_num   = 0;

    // =========================================================================
    // UART send task: bit-bang one byte LSB-first (clock-based timing)
    // =========================================================================
    task uart_send;
        input [7:0] data;
        integer i;
        begin
            @(posedge clk); #1;
            uart_rx_pin = 1'b0;  // start bit
            repeat(BAUD_CLKS) @(posedge clk);
            for (i = 0; i < 8; i = i + 1) begin
                #1;
                uart_rx_pin = data[i];
                repeat(BAUD_CLKS) @(posedge clk);
            end
            #1;
            uart_rx_pin = 1'b1;  // stop bit
            repeat(BAUD_CLKS) @(posedge clk);
        end
    endtask

    // =========================================================================
    // Helper: send a string
    // =========================================================================
    task send_string;
        input [8*80-1:0] str;  // up to 80 chars
        input integer len;
        integer i;
        reg [7:0] ch;
        begin
            for (i = 0; i < len; i = i + 1) begin
                ch = str >> ((len - 1 - i) * 8);
                uart_send(ch[7:0]);
            end
        end
    endtask

    // =========================================================================
    // Helper: send command with CR, expect OK\r\n
    // =========================================================================
    task send_command;
        input [8*20-1:0] cmd;
        input integer len;
        reg [7:0] r0, r1, r2, r3;
        begin
            send_string(cmd, len);
            uart_send(8'h0D);  // CR
            // Expect "OK\r\n"
            get_byte(r0);
            get_byte(r1);
            get_byte(r2);
            get_byte(r3);
            if (r0 !== "O" || r1 !== "K" || r2 !== 8'h0D || r3 !== 8'h0A) begin
                $display("  ERROR: expected OK\\r\\n, got 0x%02X 0x%02X 0x%02X 0x%02X",
                         r0, r1, r2, r3);
            end
        end
    endtask

    // =========================================================================
    // Helper: send command with CR, expect ERR\r\n
    // =========================================================================
    task send_command_expect_err;
        input [8*20-1:0] cmd;
        input integer len;
        reg [7:0] r0, r1, r2, r3, r4;
        begin
            send_string(cmd, len);
            uart_send(8'h0D);  // CR
            // Expect "ERR\r\n"
            get_byte(r0);
            get_byte(r1);
            get_byte(r2);
            get_byte(r3);
            get_byte(r4);
            if (r0 !== "E" || r1 !== "R" || r2 !== "R" || r3 !== 8'h0D || r4 !== 8'h0A) begin
                $display("  ERROR: expected ERR\\r\\n, got 0x%02X 0x%02X 0x%02X 0x%02X 0x%02X",
                         r0, r1, r2, r3, r4);
            end
        end
    endtask

    // =========================================================================
    // Helper: encipher a single character and return result
    // =========================================================================
    task encipher_char;
        input [7:0] pt;
        output [7:0] ct;
        begin
            uart_send(pt);
            get_byte(ct);
        end
    endtask

    // =========================================================================
    // Helper: encipher a string and check output
    // =========================================================================
    task encipher_and_check;
        input [8*40-1:0] plaintext;
        input integer pt_len;
        input [8*40-1:0] expected_ct;
        input [8*40-1:0] label;
        integer i;
        reg [7:0] pt_ch, ct_ch, exp_ch;
        reg ok;
        begin
            ok = 1'b1;
            for (i = 0; i < pt_len; i = i + 1) begin
                pt_ch = plaintext >> ((pt_len - 1 - i) * 8);
                uart_send(pt_ch[7:0]);
                get_byte(ct_ch);
                exp_ch = expected_ct >> ((pt_len - 1 - i) * 8);
                if (ct_ch !== exp_ch[7:0]) begin
                    $display("  MISMATCH at char %0d: sent '%c', expected '%c' got '%c' (0x%02X)",
                             i, pt_ch[7:0], exp_ch[7:0], ct_ch, ct_ch);
                    ok = 1'b0;
                end
            end
            if (ok) begin
                $display("PASS: %0s", label);
                pass_count = pass_count + 1;
            end else begin
                $display("FAIL: %0s", label);
                fail_count = fail_count + 1;
            end
        end
    endtask

    // =========================================================================
    // Helper: send zero-arg command (e.g. ":G", ":F", ":?")
    // These execute immediately on the opcode byte — no CR needed
    // =========================================================================
    task send_zero_arg_cmd;
        input [7:0] opcode;
        begin
            uart_send(":"); // 0x3A
            uart_send(opcode);
        end
    endtask

    // =========================================================================
    // Helper: wait for and consume banner "ENIGMA I READY\r\n"
    // =========================================================================
    task wait_for_banner;
        reg [7:0] ch;
        integer i;
        begin
            for (i = 0; i < 14; i = i + 1) begin
                get_byte(ch);
            end
            // CR
            get_byte(ch);
            if (ch !== 8'h0D) $display("  WARNING: expected CR in banner, got 0x%02X", ch);
            // LF
            get_byte(ch);
            if (ch !== 8'h0A) $display("  WARNING: expected LF in banner, got 0x%02X", ch);
        end
    endtask

    // =========================================================================
    // Helper: wait for OK\r\n
    // =========================================================================
    task wait_for_ok;
        reg [7:0] r0, r1, r2, r3;
        begin
            get_byte(r0); get_byte(r1); get_byte(r2); get_byte(r3);
            if (r0 !== "O" || r1 !== "K" || r2 !== 8'h0D || r3 !== 8'h0A)
                $display("  ERROR: expected OK, got 0x%02X('%c') 0x%02X('%c') 0x%02X 0x%02X",
                         r0, r0, r1, r1, r2, r3);
        end
    endtask

    // =========================================================================
    // Helper: send :F (factory reset), consume banner + OK
    // =========================================================================
    task factory_reset;
        begin
            send_zero_arg_cmd("F");
            wait_for_banner;
            wait_for_ok;
        end
    endtask

    // =========================================================================
    // Helper: send :G (grundstellung reset), consume OK
    // =========================================================================
    task grundstellung_reset;
        begin
            send_zero_arg_cmd("G");
            wait_for_ok;
        end
    endtask

    // =========================================================================
    // Timeout watchdog
    // =========================================================================
    initial begin
        #200_000_000_000; // 200 ms
        $display("TIMEOUT: simulation exceeded 200ms");
        $display("Results: %0d passed, %0d failed (TIMEOUT)", pass_count, fail_count);
        $finish(1);
    end

    // =========================================================================
    // Main test sequence
    // =========================================================================
    initial begin
        $display("=== FPGA Enigma I Plugboard Testbench ===");
        $display("");

        // Wait for startup banner
        wait_for_banner;
        $display("Banner received OK.");
        $display("");

        // =====================================================================
        // Test Case 1: Plugboard affects cipher output
        // Use pyenigma oracle vectors for deterministic checking.
        // Ground settings: AAAAA -> BDZGO (no plugboard)
        // With AZ plug:    AAAAA -> UTZJY
        // =====================================================================
        test_num = 1;
        $display("--- Test Case 1: Plugboard affects cipher output ---");
        factory_reset;
        send_command(":SAZ", 4);
        grundstellung_reset;
        encipher_and_check("AAAAA", 5, "UTZJY", "Case 1: AZ plugboard produces UTZJY (not BDZGO)");
        $display("");

        // =====================================================================
        // Test Case 2: :S-- clears plugboard
        // Add AZ plug, clear it, verify output returns to no-plugboard baseline.
        // =====================================================================
        test_num = 2;
        $display("--- Test Case 2: :S-- clears plugboard ---");
        factory_reset;
        send_command(":SAZ", 4);
        send_command(":S--", 4);
        grundstellung_reset;
        // After clear, should match ground settings: AAAAA -> BDZGO
        encipher_and_check("AAAAA", 5, "BDZGO", "Case 2: :S-- restores identity (BDZGO)");
        $display("");

        // =====================================================================
        // Test Case 3: Re-wire after clear
        // CD plug: HELLO -> ILBCA
        // EF plug: HELLO -> IKBDA
        // =====================================================================
        test_num = 3;
        $display("--- Test Case 3: Re-wire after clear ---");
        factory_reset;
        send_command(":SCD", 4);
        grundstellung_reset;
        encipher_and_check("HELLO", 5, "ILBCA", "Case 3a: CD plugboard (HELLO->ILBCA)");

        // Clear and re-wire with EF
        send_command(":S--", 4);
        send_command(":SEF", 4);
        grundstellung_reset;
        encipher_and_check("HELLO", 5, "IKBDA", "Case 3b: EF plugboard (HELLO->IKBDA)");
        $display("");

        // =====================================================================
        // Test Case 4: Re-wire previously wired letter after clear
        // =====================================================================
        test_num = 4;
        $display("--- Test Case 4: Re-wire previously wired letter after clear ---");

        // Add pair AB
        factory_reset;
        send_command(":SAB", 4);
        $display("  Added AB pair OK");

        // Try to add pair AC (should fail - A already wired)
        send_command_expect_err(":SAC", 4);
        $display("  AC pair rejected (A already wired) - correct");

        // Clear plugboard
        send_command(":S--", 4);
        $display("  Cleared plugboard with :S--");

        // Now AC should succeed
        send_command(":SAC", 4);
        $display("PASS: Case 4: AC pair accepted after clear (A is now free)");
        pass_count = pass_count + 1;
        $display("");

        // =====================================================================
        // Summary
        // =====================================================================
        $display("=================================");
        $display("Results: %0d passed, %0d failed", pass_count, fail_count);
        $display("=================================");
        if (fail_count == 0)
            $finish(0);
        else
            $finish(1);
    end

endmodule
